// ====================================================
/*
Project:     transactor
Engg Name:   johnson amalraj
File name:   master.sv
Description: this is the master file for transactor model
TODO :       Need to add the template
*/
// ====================================================