// ====================================================
/*
Project:     transactor
Engg Name:   johnson amalraj
File name:   env.sv
Description: this is the env file for transactor model
TODO :       Need to add the initate the master and slave
*/
// ====================================================