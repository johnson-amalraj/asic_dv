.
├── README.md
├── agenda.md
├── eda
│   ├── README.md
│   ├── default_rd_test.sv
│   ├── design.sv
│   ├── driver.sv
│   ├── env.sv
│   ├── generator.sv
│   ├── interface.sv
│   ├── random_test.sv
│   ├── tb_top.sv
│   ├── transaction.sv
│   └── wr_rd_test.sv
├── examples
│   ├── apb
│   │   ├── README.md
│   │   ├── apb_mem.sv
│   │   ├── docs
│   │   │   └── ARM_AMBA3_APB.pdf
│   │   ├── driver.sv
│   │   ├── environment.sv
│   │   ├── generator.sv
│   │   ├── interface.sv
│   │   ├── ip_monitor.sv
│   │   ├── op_monitor.sv
│   │   ├── ref_model.sv
│   │   ├── run_do.sv
│   │   ├── scoreboard.sv
│   │   ├── tb_top.sv
│   │   ├── test.sv
│   │   └── transaction.sv
│   ├── axi
│   │   ├── LICENSE
│   │   ├── README.md
│   │   ├── axi_config_objs.svh
│   │   ├── axi_env.sv
│   │   ├── axi_interface.sv
│   │   ├── axi_m_driver.sv
│   │   ├── axi_m_monitor.sv
│   │   ├── axi_master.sv
│   │   ├── axi_package.svh
│   │   ├── axi_read_seq.sv
│   │   ├── axi_s_driver.sv
│   │   ├── axi_s_monitor.sv
│   │   ├── axi_scoreboard.sv
│   │   ├── axi_slave.sv
│   │   ├── axi_tb_top.sv
│   │   ├── axi_test.sv
│   │   ├── axi_transaction.sv
│   │   ├── axi_write_seq.sv
│   │   └── docs
│   │       ├── AMBA AXI4 Specification.pdf
│   │       └── AXI.png
│   └── burst
│       ├── README.md
│       ├── env.sv
│       ├── interface.sv
│       ├── mst_agnt.sv
│       ├── mst_drvr.sv
│       ├── slv_agnt.sv
│       ├── slv_drvr.sv
│       ├── test.sv
│       └── top.sv
├── labs
│   ├── docs
│   │   ├── ECE_jS1tDVE-48-50.pdf
│   │   └── T1-System Verilog for Verification_ A Guide to Learning the Testbench Language Features.pdf
│   ├── ex1_mux_2_1
│   │   ├── basic_test.sv
│   │   ├── design.sv
│   │   ├── driver.sv
│   │   ├── environment.sv
│   │   ├── ex1_mux_2_1.sv
│   │   ├── generator.sv
│   │   ├── interface.sv
│   │   ├── testbench.sv
│   │   └── transaction.sv
│   ├── ex2_mailbox
│   │   ├── mail.sv
│   │   └── mailbox_mem.sv
│   ├── ex3_semaphore
│   │   ├── sem.sv
│   │   └── semaphore.sv
│   └── ex4_scoreboard
│       ├── default_rd_test.sv
│       ├── design.sv
│       ├── driver.sv
│       ├── environment.sv
│       ├── ex4_scoreboard.sv
│       ├── generator.sv
│       ├── interface.sv
│       ├── monitor.sv
│       ├── random_test.sv
│       ├── scoreboard.sv
│       ├── testbench.sv
│       ├── transaction.sv
│       └── wr_rd_test.sv
└── tree.sv

14 directories, 86 files
