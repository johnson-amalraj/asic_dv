// ====================================================
/*
Project:     transactor
Engg Name:   johnson amalraj
File name:   checker.sv
Description: this is the checker file for transactor model
TODO :       Need to add the template
*/
// ====================================================