// ====================================================
/*
Project:     transactor
Engg Name:   johnson amalraj
File name:   defines.sv
Description: this is the defines file for transactor model
TODO :       Need to add the required defines
*/
// ====================================================
`define HIGH = 1;
`define LOW  = 0;