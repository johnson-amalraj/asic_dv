// ====================================================
/*
Project:     transactor
Engg Name:   johnson amalraj
File name:   slave.sv
Description: this is the slave file for transactor model
TODO :       Need to add the template
*/
// ====================================================