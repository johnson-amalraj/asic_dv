// ====================================================
/*
Project:     transactor
Engg Name:   johnson amalraj
File name:   config.sv
Description: this is the config file for transactor model
TODO :       Need to add the required config
*/
// ====================================================