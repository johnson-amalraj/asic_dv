// ====================================================
/*
Project:     transactor
Engg Name:   johnson amalraj
File name:   interface.sv
Description: this is the interface file for transactor model
TODO :       Need to declare the required interface signals
*/
// ====================================================