// This is env file