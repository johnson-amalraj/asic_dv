// ====================================================
/*
Project:     transactor
Engg Name:   johnson amalraj
File name:   reg_mode.sv
Description: this is the register model file for transactor model
TODO :       Need to add the required registers
*/
// ====================================================