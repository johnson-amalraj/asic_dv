// 22-Sep-2023
