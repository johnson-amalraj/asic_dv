// ====================================================
/*
Project:     transactor
Engg Name:   johnson amalraj
File name:   asic_basic_test.sv
Description: test case for basic transaction
TODO :       Need to develop the test case
*/
// ====================================================
task asic_basic_test ();
    
endtask // endtask for asic_basic_test