// ====================================================
/*
Project:     transactor
Engg Name:   johnson amalraj
File name:   test.sv
Description: this is the test file for transactor model
TODO :       Need to connect the top and testbench
*/
// ====================================================