////////////////////////////////////////////////////////////////////////////////////////////////
// 1. Write a constraint for 8bit variables, that only give multiples of 4
////////////////////////////////////////////////////////////////////////////////////////////////

val_8b = 0;

// 0  | 00000000
// 4  | 00000100
// 8  | 00001000
// 12 | 00001100
// 16 | 00010000

// Hint : Only last 2 bits is 0, then its multiples of 4 only

constraint mul_4 {val_8b[1:0] != 0; }

////////////////////////////////////////////////////////////////////////////////////////////////
// 2. Find a clk signal frequency in time
////////////////////////////////////////////////////////////////////////////////////////////////
clk 
clk_period 

assert detect_period (clk_en)
{
disable (clk_en = 0)
(@posedge clk) ((t[0]=$realtime) -> ((@posedge clk) (t[1]=$realtime)) #0 (clk_peiod t[1]-t[0])
}

////////////////////////////////////////////////////////////////////////////////////////////////
// 3. What is inside the uvm_driver 
////////////////////////////////////////////////////////////////////////////////////////////////
main_phase()

// transaction from the sequencer

seqr.get_next_item(trans_o);
vif <= trans.addr;
vif <= trans.data;
seqr.item_done();

vrtual interface in driver

////////////////////////////////////////////////////////////////////////////////////////////////
// 4. what connection actual interface
////////////////////////////////////////////////////////////////////////////////////////////////
virtual interface VIP / normal interface DUT

////////////////////////////////////////////////////////////////////////////////////////////////
// 5. Explain uvm_env
////////////////////////////////////////////////////////////////////////////////////////////////
dut 
top
clock generation
waveform genr

dut instance (input and output)

sram

vip instance  (input output)

sram

test

env

active / passive

agent
   driver
   monitor
   sequencer

virtual interfafce 

virtual seqr.();

vritual sequencer

////////////////////////////////////////////////////////////////////////////////////////////////
// 6. out of order transactions
////////////////////////////////////////////////////////////////////////////////////////////////
scoreboard


0, 1, 2, 3
2, 4, 3

APB

DDR
addr 4, 8, 20
read 8, 4, 20

FIFO 

dynamic array
static array
assoc array

tx_arr[]
rx_arr[]

////////////////////////////////////////////////////////////////////////////////////////////////
// 7. Write a coverage for the 8bit variable, which will have only 1 in the variable
// other bins illegal bins 
////////////////////////////////////////////////////////////////////////////////////////////////

val_8b;

// onehot

valid bits 00000001
valid bits 00000010
valid bits 00000100
valid bits 00001000

coverpoint onehot_cp val_8b
{
bins 00000001 
bins 00000010 
// illegal bins 
}

function num_one (val_8b);

   if (val_8b == 1 || val_8b == 2 || val_8b = 4) begin
   end

endfunction

////////////////////////////////////////////////////////////////////////////////////////////////
// 8. scope resolution operator, what all are the places we can use it 
////////////////////////////////////////////////////////////////////////////////////////////////
import uvm_pkg::*

extern class / function :: package

////////////////////////////////////////////////////////////////////////////////////////////////
// 9. What is the difference between analysis import, export and port 
////////////////////////////////////////////////////////////////////////////////////////////////
analysis import and export

analysis_imp ()
analysis_exp

componentA

compB, compC


////////////////////////////////////////////////////////////////////////////////////////////////
// 10. How to override the soft constaint 
////////////////////////////////////////////////////////////////////////////////////////////////
rand class
constraint {;}

rand.const1

parent class

constraint A;

child class extend parent
constraint A; // should be same name as parent class
